module MEM_WB(
	input clk, 
	input rst
	);



endmodule