module WDT(
	input clk,
	input rst,
	input clk2,
	input rst2,
	input [31:0] w_addr,
	output logic WTO
	);


logic WDEN;
logic WDLIVE;
logic WTOCNT;
logic WTO;


endmodule