module CPU();


endmodule