`define Rtype 7'b0110011